`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/31/2023 02:59:56 PM
// Design Name: 
// Module Name: Register_Bank
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Register_Bank(
    input Clk,
    input [2:0] Reg_En,
    input [3:0] ValStore,
    output [3:0] Reg_0_out,
    output [3:0] Reg_1_out,
    output [3:0] Reg_2_out,
    output [3:0] Reg_3_out,
    output [3:0] Reg_4_out,
    output [3:0] Reg_5_out,
    output [3:0] Reg_6_out,
    output [3:0] Reg_7_out
    );
endmodule
